module AudPlayer(
	input i_rst_n,
	input i_bclk,
	input i_daclrck,
	input i_en, // enable AudPlayer only when playing audio, work with AudDSP
	input i_dac_data, //dac_data
	output o_aud_dacdat
);


endmodule