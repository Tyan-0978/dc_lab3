// ----------------------------------------------------------------------
// interpolation calculation module
// ----------------------------------------------------------------------

module itp5 (
    input  [15:0] i_data_1,
    input  [15:0] i_data_2,
    output [15:0] o_data_1,
    output [15:0] o_data_2,
    output [15:0] o_data_3,
    output [15:0] o_data_4,
);

endmodule

module itp6 (
    input  [15:0] i_data_1,
    input  [15:0] i_data_2,
    output [15:0] o_data_1,
    output [15:0] o_data_2,
    output [15:0] o_data_3,
    output [15:0] o_data_4,
    output [15:0] o_data_5,
);

endmodule

module itp7 (
    input  [15:0] i_data_1,
    input  [15:0] i_data_2,
    output [15:0] o_data_1,
    output [15:0] o_data_2,
    output [15:0] o_data_3,
    output [15:0] o_data_4,
    output [15:0] o_data_5,
    output [15:0] o_data_6,
);

endmodule

module itp8 (
    input  [15:0] i_data_1,
    input  [15:0] i_data_2,
    output [15:0] o_data_1,
    output [15:0] o_data_2,
    output [15:0] o_data_3,
    output [15:0] o_data_4,
    output [15:0] o_data_5,
    output [15:0] o_data_6,
    output [15:0] o_data_7,
);

endmodule
