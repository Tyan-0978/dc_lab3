// ----------------------------------------------------------------------                            
// interpolation module for slow speed
// ----------------------------------------------------------------------

module Interp (
    input         i_rst_n,
    input         i_clk,
    input         i_valid,
    input [15:0]  i_data,
    input         i_mode,
    input [3:0]   i_speed,
    output [15:0] o_slow_data,
    output        o_fetch_data
);

// ----------------------------------------------------------------------                            
// signals
// ----------------------------------------------------------------------

reg  [15:0] data_1, next_data_1;
reg  [15:0] data_2, next_data_2;

// ----------------------------------------------------------------------                            
// conbinational part
// ----------------------------------------------------------------------

// ----------------------------------------------------------------------                            
// sequential part
// ----------------------------------------------------------------------

endmodule
